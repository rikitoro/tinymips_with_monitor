// monitor.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module monitor (
		input  wire        clk_clk,            //         clk.clk
		output wire [31:0] dmem_addr_export,   //   dmem_addr.export
		output wire        dmem_clk_export,    //    dmem_clk.export
		input  wire [31:0] dmem_rd_export,     //     dmem_rd.export
		output wire [31:0] dmem_wd_export,     //     dmem_wd.export
		output wire        dmem_we_export,     //     dmem_we.export
		output wire [31:0] imem_addr_export,   //   imem_addr.export
		output wire        imem_clk_export,    //    imem_clk.export
		input  wire [31:0] imem_rd_export,     //     imem_rd.export
		output wire [31:0] imem_wd_export,     //     imem_wd.export
		output wire        imem_we_export,     //     imem_we.export
		output wire [31:0] iport3_data_export, // iport3_data.export
		input  wire [31:0] oport3_data_export, // oport3_data.export
		output wire        prg_mode_export,    //    prg_mode.export
		input  wire        reset_reset_n,      //       reset.reset_n
		output wire        rst_export,         //         rst.export
		input  wire        uart_rxd,           //        uart.rxd
		output wire        uart_txd            //            .txd
	);

	wire  [31:0] nios2_processor_data_master_readdata;                          // mm_interconnect_0:nios2_processor_data_master_readdata -> nios2_processor:d_readdata
	wire         nios2_processor_data_master_waitrequest;                       // mm_interconnect_0:nios2_processor_data_master_waitrequest -> nios2_processor:d_waitrequest
	wire         nios2_processor_data_master_debugaccess;                       // nios2_processor:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_processor_data_master_debugaccess
	wire  [15:0] nios2_processor_data_master_address;                           // nios2_processor:d_address -> mm_interconnect_0:nios2_processor_data_master_address
	wire   [3:0] nios2_processor_data_master_byteenable;                        // nios2_processor:d_byteenable -> mm_interconnect_0:nios2_processor_data_master_byteenable
	wire         nios2_processor_data_master_read;                              // nios2_processor:d_read -> mm_interconnect_0:nios2_processor_data_master_read
	wire         nios2_processor_data_master_write;                             // nios2_processor:d_write -> mm_interconnect_0:nios2_processor_data_master_write
	wire  [31:0] nios2_processor_data_master_writedata;                         // nios2_processor:d_writedata -> mm_interconnect_0:nios2_processor_data_master_writedata
	wire  [31:0] nios2_processor_instruction_master_readdata;                   // mm_interconnect_0:nios2_processor_instruction_master_readdata -> nios2_processor:i_readdata
	wire         nios2_processor_instruction_master_waitrequest;                // mm_interconnect_0:nios2_processor_instruction_master_waitrequest -> nios2_processor:i_waitrequest
	wire  [15:0] nios2_processor_instruction_master_address;                    // nios2_processor:i_address -> mm_interconnect_0:nios2_processor_instruction_master_address
	wire         nios2_processor_instruction_master_read;                       // nios2_processor:i_read -> mm_interconnect_0:nios2_processor_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;    // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;      // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;   // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;          // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;         // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;         // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;          // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios2_processor_debug_mem_slave_readdata;    // nios2_processor:debug_mem_slave_readdata -> mm_interconnect_0:nios2_processor_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_processor_debug_mem_slave_waitrequest; // nios2_processor:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_processor_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_processor_debug_mem_slave_debugaccess; // mm_interconnect_0:nios2_processor_debug_mem_slave_debugaccess -> nios2_processor:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_processor_debug_mem_slave_address;     // mm_interconnect_0:nios2_processor_debug_mem_slave_address -> nios2_processor:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_processor_debug_mem_slave_read;        // mm_interconnect_0:nios2_processor_debug_mem_slave_read -> nios2_processor:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_processor_debug_mem_slave_byteenable;  // mm_interconnect_0:nios2_processor_debug_mem_slave_byteenable -> nios2_processor:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_processor_debug_mem_slave_write;       // mm_interconnect_0:nios2_processor_debug_mem_slave_write -> nios2_processor:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_processor_debug_mem_slave_writedata;   // mm_interconnect_0:nios2_processor_debug_mem_slave_writedata -> nios2_processor:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;                 // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;                   // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire  [10:0] mm_interconnect_0_onchip_memory_s1_address;                    // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;                 // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire         mm_interconnect_0_onchip_memory_s1_write;                      // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;                  // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire         mm_interconnect_0_onchip_memory_s1_clken;                      // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire         mm_interconnect_0_imem_clk_s1_chipselect;                      // mm_interconnect_0:imem_clk_s1_chipselect -> imem_clk:chipselect
	wire  [31:0] mm_interconnect_0_imem_clk_s1_readdata;                        // imem_clk:readdata -> mm_interconnect_0:imem_clk_s1_readdata
	wire   [1:0] mm_interconnect_0_imem_clk_s1_address;                         // mm_interconnect_0:imem_clk_s1_address -> imem_clk:address
	wire         mm_interconnect_0_imem_clk_s1_write;                           // mm_interconnect_0:imem_clk_s1_write -> imem_clk:write_n
	wire  [31:0] mm_interconnect_0_imem_clk_s1_writedata;                       // mm_interconnect_0:imem_clk_s1_writedata -> imem_clk:writedata
	wire         mm_interconnect_0_imem_addr_s1_chipselect;                     // mm_interconnect_0:imem_addr_s1_chipselect -> imem_addr:chipselect
	wire  [31:0] mm_interconnect_0_imem_addr_s1_readdata;                       // imem_addr:readdata -> mm_interconnect_0:imem_addr_s1_readdata
	wire   [1:0] mm_interconnect_0_imem_addr_s1_address;                        // mm_interconnect_0:imem_addr_s1_address -> imem_addr:address
	wire         mm_interconnect_0_imem_addr_s1_write;                          // mm_interconnect_0:imem_addr_s1_write -> imem_addr:write_n
	wire  [31:0] mm_interconnect_0_imem_addr_s1_writedata;                      // mm_interconnect_0:imem_addr_s1_writedata -> imem_addr:writedata
	wire  [31:0] mm_interconnect_0_imem_rd_s1_readdata;                         // imem_rd:readdata -> mm_interconnect_0:imem_rd_s1_readdata
	wire   [1:0] mm_interconnect_0_imem_rd_s1_address;                          // mm_interconnect_0:imem_rd_s1_address -> imem_rd:address
	wire         mm_interconnect_0_imem_wd_s1_chipselect;                       // mm_interconnect_0:imem_wd_s1_chipselect -> imem_wd:chipselect
	wire  [31:0] mm_interconnect_0_imem_wd_s1_readdata;                         // imem_wd:readdata -> mm_interconnect_0:imem_wd_s1_readdata
	wire   [1:0] mm_interconnect_0_imem_wd_s1_address;                          // mm_interconnect_0:imem_wd_s1_address -> imem_wd:address
	wire         mm_interconnect_0_imem_wd_s1_write;                            // mm_interconnect_0:imem_wd_s1_write -> imem_wd:write_n
	wire  [31:0] mm_interconnect_0_imem_wd_s1_writedata;                        // mm_interconnect_0:imem_wd_s1_writedata -> imem_wd:writedata
	wire         mm_interconnect_0_dmem_we_s1_chipselect;                       // mm_interconnect_0:dmem_we_s1_chipselect -> dmem_we:chipselect
	wire  [31:0] mm_interconnect_0_dmem_we_s1_readdata;                         // dmem_we:readdata -> mm_interconnect_0:dmem_we_s1_readdata
	wire   [1:0] mm_interconnect_0_dmem_we_s1_address;                          // mm_interconnect_0:dmem_we_s1_address -> dmem_we:address
	wire         mm_interconnect_0_dmem_we_s1_write;                            // mm_interconnect_0:dmem_we_s1_write -> dmem_we:write_n
	wire  [31:0] mm_interconnect_0_dmem_we_s1_writedata;                        // mm_interconnect_0:dmem_we_s1_writedata -> dmem_we:writedata
	wire         mm_interconnect_0_dmem_addr_s1_chipselect;                     // mm_interconnect_0:dmem_addr_s1_chipselect -> dmem_addr:chipselect
	wire  [31:0] mm_interconnect_0_dmem_addr_s1_readdata;                       // dmem_addr:readdata -> mm_interconnect_0:dmem_addr_s1_readdata
	wire   [1:0] mm_interconnect_0_dmem_addr_s1_address;                        // mm_interconnect_0:dmem_addr_s1_address -> dmem_addr:address
	wire         mm_interconnect_0_dmem_addr_s1_write;                          // mm_interconnect_0:dmem_addr_s1_write -> dmem_addr:write_n
	wire  [31:0] mm_interconnect_0_dmem_addr_s1_writedata;                      // mm_interconnect_0:dmem_addr_s1_writedata -> dmem_addr:writedata
	wire  [31:0] mm_interconnect_0_dmem_rd_s1_readdata;                         // dmem_rd:readdata -> mm_interconnect_0:dmem_rd_s1_readdata
	wire   [1:0] mm_interconnect_0_dmem_rd_s1_address;                          // mm_interconnect_0:dmem_rd_s1_address -> dmem_rd:address
	wire         mm_interconnect_0_dmem_wd_s1_chipselect;                       // mm_interconnect_0:dmem_wd_s1_chipselect -> dmem_wd:chipselect
	wire  [31:0] mm_interconnect_0_dmem_wd_s1_readdata;                         // dmem_wd:readdata -> mm_interconnect_0:dmem_wd_s1_readdata
	wire   [1:0] mm_interconnect_0_dmem_wd_s1_address;                          // mm_interconnect_0:dmem_wd_s1_address -> dmem_wd:address
	wire         mm_interconnect_0_dmem_wd_s1_write;                            // mm_interconnect_0:dmem_wd_s1_write -> dmem_wd:write_n
	wire  [31:0] mm_interconnect_0_dmem_wd_s1_writedata;                        // mm_interconnect_0:dmem_wd_s1_writedata -> dmem_wd:writedata
	wire         mm_interconnect_0_prg_mode_s1_chipselect;                      // mm_interconnect_0:prg_mode_s1_chipselect -> prg_mode:chipselect
	wire  [31:0] mm_interconnect_0_prg_mode_s1_readdata;                        // prg_mode:readdata -> mm_interconnect_0:prg_mode_s1_readdata
	wire   [1:0] mm_interconnect_0_prg_mode_s1_address;                         // mm_interconnect_0:prg_mode_s1_address -> prg_mode:address
	wire         mm_interconnect_0_prg_mode_s1_write;                           // mm_interconnect_0:prg_mode_s1_write -> prg_mode:write_n
	wire  [31:0] mm_interconnect_0_prg_mode_s1_writedata;                       // mm_interconnect_0:prg_mode_s1_writedata -> prg_mode:writedata
	wire         mm_interconnect_0_rst_s1_chipselect;                           // mm_interconnect_0:rst_s1_chipselect -> rst:chipselect
	wire  [31:0] mm_interconnect_0_rst_s1_readdata;                             // rst:readdata -> mm_interconnect_0:rst_s1_readdata
	wire   [1:0] mm_interconnect_0_rst_s1_address;                              // mm_interconnect_0:rst_s1_address -> rst:address
	wire         mm_interconnect_0_rst_s1_write;                                // mm_interconnect_0:rst_s1_write -> rst:write_n
	wire  [31:0] mm_interconnect_0_rst_s1_writedata;                            // mm_interconnect_0:rst_s1_writedata -> rst:writedata
	wire         mm_interconnect_0_iport3_data_s1_chipselect;                   // mm_interconnect_0:iport3_data_s1_chipselect -> iport3_data:chipselect
	wire  [31:0] mm_interconnect_0_iport3_data_s1_readdata;                     // iport3_data:readdata -> mm_interconnect_0:iport3_data_s1_readdata
	wire   [1:0] mm_interconnect_0_iport3_data_s1_address;                      // mm_interconnect_0:iport3_data_s1_address -> iport3_data:address
	wire         mm_interconnect_0_iport3_data_s1_write;                        // mm_interconnect_0:iport3_data_s1_write -> iport3_data:write_n
	wire  [31:0] mm_interconnect_0_iport3_data_s1_writedata;                    // mm_interconnect_0:iport3_data_s1_writedata -> iport3_data:writedata
	wire  [31:0] mm_interconnect_0_oport3_data_s1_readdata;                     // oport3_data:readdata -> mm_interconnect_0:oport3_data_s1_readdata
	wire   [1:0] mm_interconnect_0_oport3_data_s1_address;                      // mm_interconnect_0:oport3_data_s1_address -> oport3_data:address
	wire         mm_interconnect_0_uart_s1_chipselect;                          // mm_interconnect_0:uart_s1_chipselect -> uart:chipselect
	wire  [15:0] mm_interconnect_0_uart_s1_readdata;                            // uart:readdata -> mm_interconnect_0:uart_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_s1_address;                             // mm_interconnect_0:uart_s1_address -> uart:address
	wire         mm_interconnect_0_uart_s1_read;                                // mm_interconnect_0:uart_s1_read -> uart:read_n
	wire         mm_interconnect_0_uart_s1_begintransfer;                       // mm_interconnect_0:uart_s1_begintransfer -> uart:begintransfer
	wire         mm_interconnect_0_uart_s1_write;                               // mm_interconnect_0:uart_s1_write -> uart:write_n
	wire  [15:0] mm_interconnect_0_uart_s1_writedata;                           // mm_interconnect_0:uart_s1_writedata -> uart:writedata
	wire         mm_interconnect_0_imem_we_s1_chipselect;                       // mm_interconnect_0:imem_we_s1_chipselect -> imem_we:chipselect
	wire  [31:0] mm_interconnect_0_imem_we_s1_readdata;                         // imem_we:readdata -> mm_interconnect_0:imem_we_s1_readdata
	wire   [1:0] mm_interconnect_0_imem_we_s1_address;                          // mm_interconnect_0:imem_we_s1_address -> imem_we:address
	wire         mm_interconnect_0_imem_we_s1_write;                            // mm_interconnect_0:imem_we_s1_write -> imem_we:write_n
	wire  [31:0] mm_interconnect_0_imem_we_s1_writedata;                        // mm_interconnect_0:imem_we_s1_writedata -> imem_we:writedata
	wire         mm_interconnect_0_dmem_clk_s1_chipselect;                      // mm_interconnect_0:dmem_clk_s1_chipselect -> dmem_clk:chipselect
	wire  [31:0] mm_interconnect_0_dmem_clk_s1_readdata;                        // dmem_clk:readdata -> mm_interconnect_0:dmem_clk_s1_readdata
	wire   [1:0] mm_interconnect_0_dmem_clk_s1_address;                         // mm_interconnect_0:dmem_clk_s1_address -> dmem_clk:address
	wire         mm_interconnect_0_dmem_clk_s1_write;                           // mm_interconnect_0:dmem_clk_s1_write -> dmem_clk:write_n
	wire  [31:0] mm_interconnect_0_dmem_clk_s1_writedata;                       // mm_interconnect_0:dmem_clk_s1_writedata -> dmem_clk:writedata
	wire         irq_mapper_receiver0_irq;                                      // uart:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                      // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_processor_irq_irq;                                       // irq_mapper:sender_irq -> nios2_processor:irq
	wire         rst_controller_reset_out_reset;                                // rst_controller:reset_out -> [dmem_addr:reset_n, dmem_clk:reset_n, dmem_rd:reset_n, dmem_wd:reset_n, dmem_we:reset_n, imem_addr:reset_n, imem_clk:reset_n, imem_rd:reset_n, imem_wd:reset_n, imem_we:reset_n, iport3_data:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_processor_reset_reset_bridge_in_reset_reset, nios2_processor:reset_n, onchip_memory:reset, oport3_data:reset_n, prg_mode:reset_n, rst:reset_n, rst_translator:in_reset, sysid_qsys_0:reset_n, uart:reset_n]
	wire         rst_controller_reset_out_reset_req;                            // rst_controller:reset_req -> [nios2_processor:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]

	monitor_dmem_addr dmem_addr (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_dmem_addr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dmem_addr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dmem_addr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dmem_addr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dmem_addr_s1_readdata),   //                    .readdata
		.out_port   (dmem_addr_export)                           // external_connection.export
	);

	monitor_dmem_clk dmem_clk (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_dmem_clk_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dmem_clk_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dmem_clk_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dmem_clk_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dmem_clk_s1_readdata),   //                    .readdata
		.out_port   (dmem_clk_export)                           // external_connection.export
	);

	monitor_dmem_rd dmem_rd (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_dmem_rd_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_dmem_rd_s1_readdata), //                    .readdata
		.in_port  (dmem_rd_export)                         // external_connection.export
	);

	monitor_dmem_addr dmem_wd (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_dmem_wd_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dmem_wd_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dmem_wd_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dmem_wd_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dmem_wd_s1_readdata),   //                    .readdata
		.out_port   (dmem_wd_export)                           // external_connection.export
	);

	monitor_dmem_clk dmem_we (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_dmem_we_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dmem_we_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dmem_we_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dmem_we_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dmem_we_s1_readdata),   //                    .readdata
		.out_port   (dmem_we_export)                           // external_connection.export
	);

	monitor_dmem_addr imem_addr (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_imem_addr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_imem_addr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_imem_addr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_imem_addr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_imem_addr_s1_readdata),   //                    .readdata
		.out_port   (imem_addr_export)                           // external_connection.export
	);

	monitor_dmem_clk imem_clk (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_imem_clk_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_imem_clk_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_imem_clk_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_imem_clk_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_imem_clk_s1_readdata),   //                    .readdata
		.out_port   (imem_clk_export)                           // external_connection.export
	);

	monitor_dmem_rd imem_rd (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_imem_rd_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_imem_rd_s1_readdata), //                    .readdata
		.in_port  (imem_rd_export)                         // external_connection.export
	);

	monitor_dmem_addr imem_wd (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_imem_wd_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_imem_wd_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_imem_wd_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_imem_wd_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_imem_wd_s1_readdata),   //                    .readdata
		.out_port   (imem_wd_export)                           // external_connection.export
	);

	monitor_dmem_clk imem_we (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_imem_we_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_imem_we_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_imem_we_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_imem_we_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_imem_we_s1_readdata),   //                    .readdata
		.out_port   (imem_we_export)                           // external_connection.export
	);

	monitor_dmem_addr iport3_data (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_iport3_data_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_iport3_data_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_iport3_data_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_iport3_data_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_iport3_data_s1_readdata),   //                    .readdata
		.out_port   (iport3_data_export)                           // external_connection.export
	);

	monitor_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                     //               irq.irq
	);

	monitor_nios2_processor nios2_processor (
		.clk                                 (clk_clk),                                                       //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                               //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                            //                          .reset_req
		.d_address                           (nios2_processor_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_processor_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_processor_data_master_read),                              //                          .read
		.d_readdata                          (nios2_processor_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_processor_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_processor_data_master_write),                             //                          .write
		.d_writedata                         (nios2_processor_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_processor_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_processor_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_processor_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_processor_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_processor_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_processor_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                              //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_processor_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_processor_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_processor_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_processor_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_processor_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_processor_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_processor_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_processor_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                               // custom_instruction_master.readra
	);

	monitor_onchip_memory onchip_memory (
		.clk        (clk_clk),                                       //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)             //       .reset_req
	);

	monitor_dmem_rd oport3_data (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_oport3_data_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_oport3_data_s1_readdata), //                    .readdata
		.in_port  (oport3_data_export)                         // external_connection.export
	);

	monitor_dmem_clk prg_mode (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_prg_mode_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_prg_mode_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_prg_mode_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_prg_mode_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_prg_mode_s1_readdata),   //                    .readdata
		.out_port   (prg_mode_export)                           // external_connection.export
	);

	monitor_dmem_clk rst (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_rst_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_rst_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_rst_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_rst_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_rst_s1_readdata),   //                    .readdata
		.out_port   (rst_export)                           // external_connection.export
	);

	monitor_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	monitor_uart uart (
		.clk           (clk_clk),                                 //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address       (mm_interconnect_0_uart_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_s1_readdata),      //                    .readdata
		.dataavailable (),                                        //                    .dataavailable
		.readyfordata  (),                                        //                    .readyfordata
		.rxd           (uart_rxd),                                // external_connection.export
		.txd           (uart_txd),                                //                    .export
		.irq           (irq_mapper_receiver0_irq)                 //                 irq.irq
	);

	monitor_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                     (clk_clk),                                                       //                                   clk_0_clk.clk
		.nios2_processor_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                // nios2_processor_reset_reset_bridge_in_reset.reset
		.nios2_processor_data_master_address               (nios2_processor_data_master_address),                           //                 nios2_processor_data_master.address
		.nios2_processor_data_master_waitrequest           (nios2_processor_data_master_waitrequest),                       //                                            .waitrequest
		.nios2_processor_data_master_byteenable            (nios2_processor_data_master_byteenable),                        //                                            .byteenable
		.nios2_processor_data_master_read                  (nios2_processor_data_master_read),                              //                                            .read
		.nios2_processor_data_master_readdata              (nios2_processor_data_master_readdata),                          //                                            .readdata
		.nios2_processor_data_master_write                 (nios2_processor_data_master_write),                             //                                            .write
		.nios2_processor_data_master_writedata             (nios2_processor_data_master_writedata),                         //                                            .writedata
		.nios2_processor_data_master_debugaccess           (nios2_processor_data_master_debugaccess),                       //                                            .debugaccess
		.nios2_processor_instruction_master_address        (nios2_processor_instruction_master_address),                    //          nios2_processor_instruction_master.address
		.nios2_processor_instruction_master_waitrequest    (nios2_processor_instruction_master_waitrequest),                //                                            .waitrequest
		.nios2_processor_instruction_master_read           (nios2_processor_instruction_master_read),                       //                                            .read
		.nios2_processor_instruction_master_readdata       (nios2_processor_instruction_master_readdata),                   //                                            .readdata
		.dmem_addr_s1_address                              (mm_interconnect_0_dmem_addr_s1_address),                        //                                dmem_addr_s1.address
		.dmem_addr_s1_write                                (mm_interconnect_0_dmem_addr_s1_write),                          //                                            .write
		.dmem_addr_s1_readdata                             (mm_interconnect_0_dmem_addr_s1_readdata),                       //                                            .readdata
		.dmem_addr_s1_writedata                            (mm_interconnect_0_dmem_addr_s1_writedata),                      //                                            .writedata
		.dmem_addr_s1_chipselect                           (mm_interconnect_0_dmem_addr_s1_chipselect),                     //                                            .chipselect
		.dmem_clk_s1_address                               (mm_interconnect_0_dmem_clk_s1_address),                         //                                 dmem_clk_s1.address
		.dmem_clk_s1_write                                 (mm_interconnect_0_dmem_clk_s1_write),                           //                                            .write
		.dmem_clk_s1_readdata                              (mm_interconnect_0_dmem_clk_s1_readdata),                        //                                            .readdata
		.dmem_clk_s1_writedata                             (mm_interconnect_0_dmem_clk_s1_writedata),                       //                                            .writedata
		.dmem_clk_s1_chipselect                            (mm_interconnect_0_dmem_clk_s1_chipselect),                      //                                            .chipselect
		.dmem_rd_s1_address                                (mm_interconnect_0_dmem_rd_s1_address),                          //                                  dmem_rd_s1.address
		.dmem_rd_s1_readdata                               (mm_interconnect_0_dmem_rd_s1_readdata),                         //                                            .readdata
		.dmem_wd_s1_address                                (mm_interconnect_0_dmem_wd_s1_address),                          //                                  dmem_wd_s1.address
		.dmem_wd_s1_write                                  (mm_interconnect_0_dmem_wd_s1_write),                            //                                            .write
		.dmem_wd_s1_readdata                               (mm_interconnect_0_dmem_wd_s1_readdata),                         //                                            .readdata
		.dmem_wd_s1_writedata                              (mm_interconnect_0_dmem_wd_s1_writedata),                        //                                            .writedata
		.dmem_wd_s1_chipselect                             (mm_interconnect_0_dmem_wd_s1_chipselect),                       //                                            .chipselect
		.dmem_we_s1_address                                (mm_interconnect_0_dmem_we_s1_address),                          //                                  dmem_we_s1.address
		.dmem_we_s1_write                                  (mm_interconnect_0_dmem_we_s1_write),                            //                                            .write
		.dmem_we_s1_readdata                               (mm_interconnect_0_dmem_we_s1_readdata),                         //                                            .readdata
		.dmem_we_s1_writedata                              (mm_interconnect_0_dmem_we_s1_writedata),                        //                                            .writedata
		.dmem_we_s1_chipselect                             (mm_interconnect_0_dmem_we_s1_chipselect),                       //                                            .chipselect
		.imem_addr_s1_address                              (mm_interconnect_0_imem_addr_s1_address),                        //                                imem_addr_s1.address
		.imem_addr_s1_write                                (mm_interconnect_0_imem_addr_s1_write),                          //                                            .write
		.imem_addr_s1_readdata                             (mm_interconnect_0_imem_addr_s1_readdata),                       //                                            .readdata
		.imem_addr_s1_writedata                            (mm_interconnect_0_imem_addr_s1_writedata),                      //                                            .writedata
		.imem_addr_s1_chipselect                           (mm_interconnect_0_imem_addr_s1_chipselect),                     //                                            .chipselect
		.imem_clk_s1_address                               (mm_interconnect_0_imem_clk_s1_address),                         //                                 imem_clk_s1.address
		.imem_clk_s1_write                                 (mm_interconnect_0_imem_clk_s1_write),                           //                                            .write
		.imem_clk_s1_readdata                              (mm_interconnect_0_imem_clk_s1_readdata),                        //                                            .readdata
		.imem_clk_s1_writedata                             (mm_interconnect_0_imem_clk_s1_writedata),                       //                                            .writedata
		.imem_clk_s1_chipselect                            (mm_interconnect_0_imem_clk_s1_chipselect),                      //                                            .chipselect
		.imem_rd_s1_address                                (mm_interconnect_0_imem_rd_s1_address),                          //                                  imem_rd_s1.address
		.imem_rd_s1_readdata                               (mm_interconnect_0_imem_rd_s1_readdata),                         //                                            .readdata
		.imem_wd_s1_address                                (mm_interconnect_0_imem_wd_s1_address),                          //                                  imem_wd_s1.address
		.imem_wd_s1_write                                  (mm_interconnect_0_imem_wd_s1_write),                            //                                            .write
		.imem_wd_s1_readdata                               (mm_interconnect_0_imem_wd_s1_readdata),                         //                                            .readdata
		.imem_wd_s1_writedata                              (mm_interconnect_0_imem_wd_s1_writedata),                        //                                            .writedata
		.imem_wd_s1_chipselect                             (mm_interconnect_0_imem_wd_s1_chipselect),                       //                                            .chipselect
		.imem_we_s1_address                                (mm_interconnect_0_imem_we_s1_address),                          //                                  imem_we_s1.address
		.imem_we_s1_write                                  (mm_interconnect_0_imem_we_s1_write),                            //                                            .write
		.imem_we_s1_readdata                               (mm_interconnect_0_imem_we_s1_readdata),                         //                                            .readdata
		.imem_we_s1_writedata                              (mm_interconnect_0_imem_we_s1_writedata),                        //                                            .writedata
		.imem_we_s1_chipselect                             (mm_interconnect_0_imem_we_s1_chipselect),                       //                                            .chipselect
		.iport3_data_s1_address                            (mm_interconnect_0_iport3_data_s1_address),                      //                              iport3_data_s1.address
		.iport3_data_s1_write                              (mm_interconnect_0_iport3_data_s1_write),                        //                                            .write
		.iport3_data_s1_readdata                           (mm_interconnect_0_iport3_data_s1_readdata),                     //                                            .readdata
		.iport3_data_s1_writedata                          (mm_interconnect_0_iport3_data_s1_writedata),                    //                                            .writedata
		.iport3_data_s1_chipselect                         (mm_interconnect_0_iport3_data_s1_chipselect),                   //                                            .chipselect
		.jtag_uart_0_avalon_jtag_slave_address             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),       //               jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),         //                                            .write
		.jtag_uart_0_avalon_jtag_slave_read                (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),          //                                            .read
		.jtag_uart_0_avalon_jtag_slave_readdata            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),      //                                            .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),     //                                            .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),   //                                            .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),    //                                            .chipselect
		.nios2_processor_debug_mem_slave_address           (mm_interconnect_0_nios2_processor_debug_mem_slave_address),     //             nios2_processor_debug_mem_slave.address
		.nios2_processor_debug_mem_slave_write             (mm_interconnect_0_nios2_processor_debug_mem_slave_write),       //                                            .write
		.nios2_processor_debug_mem_slave_read              (mm_interconnect_0_nios2_processor_debug_mem_slave_read),        //                                            .read
		.nios2_processor_debug_mem_slave_readdata          (mm_interconnect_0_nios2_processor_debug_mem_slave_readdata),    //                                            .readdata
		.nios2_processor_debug_mem_slave_writedata         (mm_interconnect_0_nios2_processor_debug_mem_slave_writedata),   //                                            .writedata
		.nios2_processor_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_processor_debug_mem_slave_byteenable),  //                                            .byteenable
		.nios2_processor_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_processor_debug_mem_slave_waitrequest), //                                            .waitrequest
		.nios2_processor_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_processor_debug_mem_slave_debugaccess), //                                            .debugaccess
		.onchip_memory_s1_address                          (mm_interconnect_0_onchip_memory_s1_address),                    //                            onchip_memory_s1.address
		.onchip_memory_s1_write                            (mm_interconnect_0_onchip_memory_s1_write),                      //                                            .write
		.onchip_memory_s1_readdata                         (mm_interconnect_0_onchip_memory_s1_readdata),                   //                                            .readdata
		.onchip_memory_s1_writedata                        (mm_interconnect_0_onchip_memory_s1_writedata),                  //                                            .writedata
		.onchip_memory_s1_byteenable                       (mm_interconnect_0_onchip_memory_s1_byteenable),                 //                                            .byteenable
		.onchip_memory_s1_chipselect                       (mm_interconnect_0_onchip_memory_s1_chipselect),                 //                                            .chipselect
		.onchip_memory_s1_clken                            (mm_interconnect_0_onchip_memory_s1_clken),                      //                                            .clken
		.oport3_data_s1_address                            (mm_interconnect_0_oport3_data_s1_address),                      //                              oport3_data_s1.address
		.oport3_data_s1_readdata                           (mm_interconnect_0_oport3_data_s1_readdata),                     //                                            .readdata
		.prg_mode_s1_address                               (mm_interconnect_0_prg_mode_s1_address),                         //                                 prg_mode_s1.address
		.prg_mode_s1_write                                 (mm_interconnect_0_prg_mode_s1_write),                           //                                            .write
		.prg_mode_s1_readdata                              (mm_interconnect_0_prg_mode_s1_readdata),                        //                                            .readdata
		.prg_mode_s1_writedata                             (mm_interconnect_0_prg_mode_s1_writedata),                       //                                            .writedata
		.prg_mode_s1_chipselect                            (mm_interconnect_0_prg_mode_s1_chipselect),                      //                                            .chipselect
		.rst_s1_address                                    (mm_interconnect_0_rst_s1_address),                              //                                      rst_s1.address
		.rst_s1_write                                      (mm_interconnect_0_rst_s1_write),                                //                                            .write
		.rst_s1_readdata                                   (mm_interconnect_0_rst_s1_readdata),                             //                                            .readdata
		.rst_s1_writedata                                  (mm_interconnect_0_rst_s1_writedata),                            //                                            .writedata
		.rst_s1_chipselect                                 (mm_interconnect_0_rst_s1_chipselect),                           //                                            .chipselect
		.sysid_qsys_0_control_slave_address                (mm_interconnect_0_sysid_qsys_0_control_slave_address),          //                  sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata               (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),         //                                            .readdata
		.uart_s1_address                                   (mm_interconnect_0_uart_s1_address),                             //                                     uart_s1.address
		.uart_s1_write                                     (mm_interconnect_0_uart_s1_write),                               //                                            .write
		.uart_s1_read                                      (mm_interconnect_0_uart_s1_read),                                //                                            .read
		.uart_s1_readdata                                  (mm_interconnect_0_uart_s1_readdata),                            //                                            .readdata
		.uart_s1_writedata                                 (mm_interconnect_0_uart_s1_writedata),                           //                                            .writedata
		.uart_s1_begintransfer                             (mm_interconnect_0_uart_s1_begintransfer),                       //                                            .begintransfer
		.uart_s1_chipselect                                (mm_interconnect_0_uart_s1_chipselect)                           //                                            .chipselect
	);

	monitor_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_processor_irq_irq)         //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
